// mcu_qsys.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module mcu_qsys (
		input  wire        clk_clk,                          //               clk.clk
		output wire [66:0] hps_0_h2f_loan_io_in,             // hps_0_h2f_loan_io.in
		input  wire [66:0] hps_0_h2f_loan_io_out,            //                  .out
		input  wire [66:0] hps_0_h2f_loan_io_oe,             //                  .oe
		input  wire        hps_0_uart0_cts,                  //       hps_0_uart0.cts
		input  wire        hps_0_uart0_dsr,                  //                  .dsr
		input  wire        hps_0_uart0_dcd,                  //                  .dcd
		input  wire        hps_0_uart0_ri,                   //                  .ri
		output wire        hps_0_uart0_dtr,                  //                  .dtr
		output wire        hps_0_uart0_rts,                  //                  .rts
		output wire        hps_0_uart0_out1_n,               //                  .out1_n
		output wire        hps_0_uart0_out2_n,               //                  .out2_n
		input  wire        hps_0_uart0_rxd,                  //                  .rxd
		output wire        hps_0_uart0_txd,                  //                  .txd
		inout  wire        hps_io_hps_io_gpio_inst_LOANIO49, //            hps_io.hps_io_gpio_inst_LOANIO49
		inout  wire        hps_io_hps_io_gpio_inst_LOANIO50, //                  .hps_io_gpio_inst_LOANIO50
		output wire [12:0] memory_mem_a,                     //            memory.mem_a
		output wire [2:0]  memory_mem_ba,                    //                  .mem_ba
		output wire        memory_mem_ck,                    //                  .mem_ck
		output wire        memory_mem_ck_n,                  //                  .mem_ck_n
		output wire        memory_mem_cke,                   //                  .mem_cke
		output wire        memory_mem_cs_n,                  //                  .mem_cs_n
		output wire        memory_mem_ras_n,                 //                  .mem_ras_n
		output wire        memory_mem_cas_n,                 //                  .mem_cas_n
		output wire        memory_mem_we_n,                  //                  .mem_we_n
		output wire        memory_mem_reset_n,               //                  .mem_reset_n
		inout  wire [7:0]  memory_mem_dq,                    //                  .mem_dq
		inout  wire        memory_mem_dqs,                   //                  .mem_dqs
		inout  wire        memory_mem_dqs_n,                 //                  .mem_dqs_n
		output wire        memory_mem_odt,                   //                  .mem_odt
		output wire        memory_mem_dm,                    //                  .mem_dm
		input  wire        memory_oct_rzqin,                 //                  .oct_rzqin
		input  wire        reset_reset_n                     //             reset.reset_n
	);

	mcu_qsys_hps_0 #(
		.F2S_Width (0),
		.S2F_Width (0)
	) hps_0 (
		.h2f_loan_in               (hps_0_h2f_loan_io_in),             // h2f_loan_io.in
		.h2f_loan_out              (hps_0_h2f_loan_io_out),            //            .out
		.h2f_loan_oe               (hps_0_h2f_loan_io_oe),             //            .oe
		.uart0_cts                 (hps_0_uart0_cts),                  //       uart0.cts
		.uart0_dsr                 (hps_0_uart0_dsr),                  //            .dsr
		.uart0_dcd                 (hps_0_uart0_dcd),                  //            .dcd
		.uart0_ri                  (hps_0_uart0_ri),                   //            .ri
		.uart0_dtr                 (hps_0_uart0_dtr),                  //            .dtr
		.uart0_rts                 (hps_0_uart0_rts),                  //            .rts
		.uart0_out1_n              (hps_0_uart0_out1_n),               //            .out1_n
		.uart0_out2_n              (hps_0_uart0_out2_n),               //            .out2_n
		.uart0_rxd                 (hps_0_uart0_rxd),                  //            .rxd
		.uart0_txd                 (hps_0_uart0_txd),                  //            .txd
		.mem_a                     (memory_mem_a),                     //      memory.mem_a
		.mem_ba                    (memory_mem_ba),                    //            .mem_ba
		.mem_ck                    (memory_mem_ck),                    //            .mem_ck
		.mem_ck_n                  (memory_mem_ck_n),                  //            .mem_ck_n
		.mem_cke                   (memory_mem_cke),                   //            .mem_cke
		.mem_cs_n                  (memory_mem_cs_n),                  //            .mem_cs_n
		.mem_ras_n                 (memory_mem_ras_n),                 //            .mem_ras_n
		.mem_cas_n                 (memory_mem_cas_n),                 //            .mem_cas_n
		.mem_we_n                  (memory_mem_we_n),                  //            .mem_we_n
		.mem_reset_n               (memory_mem_reset_n),               //            .mem_reset_n
		.mem_dq                    (memory_mem_dq),                    //            .mem_dq
		.mem_dqs                   (memory_mem_dqs),                   //            .mem_dqs
		.mem_dqs_n                 (memory_mem_dqs_n),                 //            .mem_dqs_n
		.mem_odt                   (memory_mem_odt),                   //            .mem_odt
		.mem_dm                    (memory_mem_dm),                    //            .mem_dm
		.oct_rzqin                 (memory_oct_rzqin),                 //            .oct_rzqin
		.hps_io_gpio_inst_LOANIO49 (hps_io_hps_io_gpio_inst_LOANIO49), //      hps_io.hps_io_gpio_inst_LOANIO49
		.hps_io_gpio_inst_LOANIO50 (hps_io_hps_io_gpio_inst_LOANIO50), //            .hps_io_gpio_inst_LOANIO50
		.h2f_rst_n                 ()                                  //   h2f_reset.reset_n
	);

endmodule
