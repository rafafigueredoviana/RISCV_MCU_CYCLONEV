// Copyright 2017 ETH Zurich and University of Bologna.
// Copyright and related rights are licensed under the Solderpad Hardware
// License, Version 0.51 (the “License”); you may not use this file except in
// compliance with the License.  You may obtain a copy of the License at
// http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
// or agreed to in writing, software, hardware and materials distributed under
// this License is distributed on an “AS IS” BASIS, WITHOUT WARRANTIES OR
// CONDITIONS OF ANY KIND, either express or implied. See the License for the
// specific language governing permissions and limitations under the License.

`ifndef CONFIG_SV
`define CONFIG_SV
  `define RISCV
  `define SIMULATION
  // `define PULP_FPGA_EMUL
  // always define ASIC when we do a synthesis run
  `ifndef SIMULATION
    `ifndef PULP_FPGA_EMUL
      `ifdef SYNTHESIS
        `define ASIC
      `endif
    `endif
  `endif
  // data and instruction RAM address and word width
  `define ROM_ADDR_WIDTH      12
  `define ROM_START_ADDR      32'h8000

  // General defines

  `define AXI_ADDR_WIDTH       = 32,
  `define AXI_DATA_WIDTH       = 32,
  `define AXI_ID_MASTER_WIDTH  = 2,
  `define AXI_ID_SLAVE_WIDTH   = 2,
  `define AXI_USER_WIDTH       = 0,
  `define APB_ADDR_WIDTH       = 32,
  `define APB_DATA_WIDTH       = 32,
  `define DATA_RAM_SIZE        = 32768, // in bytes
  `define INSTR_RAM_SIZE       = 32768, // in bytes
  `define USE_ZERO_RISCY       = 0,
  `define RISCY_RV32F          = 1,
  `define ZERO_RV32M           = 0,
  `define ZERO_RV32E           = 0

  // Simulation only stuff
  `ifndef SYNTHESIS
  //`define DATA_STALL_RANDOM
  //`define INSTR_STALL_RANDOM
  `endif

`endif
